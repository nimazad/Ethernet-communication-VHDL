`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Create Date:    Wed May 19 17:16:14 2010
// Design Name: 
// Module Name:    netlist_1_EMPTY
//////////////////////////////////////////////////////////////////////////////////
module netlist_1_EMPTY(In_CLK_50_Ref_E1, In_PHY_RX0_J9, In_PHY_RX1_J8, In_PHY_CRS_G13, Out_PHY_DATA_0_D3, Out_PHY_DATA_1_F4, Out_PHY_TXEN_E4, Out_PHY_MDIO_J7, Out_PHY_MDC_H6, Out_PHY_Reset_J6, Out_LED_C0_AC1, Out_LED_C1_AB1, Out_LED_C2_W6, Out_RP6_AF14, Out_RP4_AD15, Out_RP8_AE14, Out_RP9_AF13, Out_RP18_P1, Out_RP17_M2, R_EXTCLK_A14, R_FRAME_VALID_F20, R_LINE_VALID_F19, R_PIXCLK_C16, R_TRIGGER_A15, R_CAM_DATA0_C22, R_CAM_DATA1_D22, R_CAM_DATA2_C23, R_CAM_DATA3_D23, R_CAM_DATA4_A22, R_CAM_DATA5_B23, R_CAM_DATA6_G17, R_CAM_DATA7_H17, R_CAM_DATA8_B21, R_CAM_DATA9_C21, R_CAM_DATA10_D21, R_CAM_DATA11_E21, L_EXTCLK_B13, L_FRAME_VALID_F12, L_LINE_VALID_C11, L_PIXCLK_K11, L_TRIGGER_G10, L_CAM_DATA0_B10, L_CAM_DATA1_A10, L_CAM_DATA2_D10, L_CAM_DATA3_C10, L_CAM_DATA4_H12, L_CAM_DATA5_G12, L_CAM_DATA6_B9, L_CAM_DATA7_A9, L_CAM_DATA8_D9, L_CAM_DATA9_E10, L_CAM_DATA10_B8, L_CAM_DATA11_C7, InOut_I2C_L_SDA_B15, InOut_I2C_L_SCL_F14, InOut_I2C_R_SDA_G9, InOut_I2C_R_SCL_F7);
  input In_CLK_50_Ref_E1;
  input In_PHY_RX0_J9;
  input In_PHY_RX1_J8;
  input In_PHY_CRS_G13;
  output Out_PHY_DATA_0_D3;
  output Out_PHY_DATA_1_F4;
  output Out_PHY_TXEN_E4;
  inout  Out_PHY_MDIO_J7;
  output Out_PHY_MDC_H6;
  output Out_PHY_Reset_J6;
  output Out_LED_C0_AC1;
  output Out_LED_C1_AB1;
  output Out_LED_C2_W6;
  output Out_RP6_AF14;
  output Out_RP4_AD15;
  output Out_RP8_AE14;
  output Out_RP9_AF13;
  output Out_RP18_P1;
  output Out_RP17_M2;
  input R_EXTCLK_A14;
  input R_FRAME_VALID_F20;
  input R_LINE_VALID_F19;
  input R_PIXCLK_C16;
  output R_TRIGGER_A15;
  input R_CAM_DATA0_C22;
  input R_CAM_DATA1_D22;
  input R_CAM_DATA2_C23;
  input R_CAM_DATA3_D23;
  input R_CAM_DATA4_A22;
  input R_CAM_DATA5_B23;
  input R_CAM_DATA6_G17;
  input R_CAM_DATA7_H17;
  input R_CAM_DATA8_B21;
  input R_CAM_DATA9_C21;
  input R_CAM_DATA10_D21;
  input R_CAM_DATA11_E21;
  input L_EXTCLK_B13;
  input L_FRAME_VALID_F12;
  input L_LINE_VALID_C11;
  input L_PIXCLK_K11;
  output L_TRIGGER_G10;
  input L_CAM_DATA0_B10;
  input L_CAM_DATA1_A10;
  input L_CAM_DATA2_D10;
  input L_CAM_DATA3_C10;
  input L_CAM_DATA4_H12;
  input L_CAM_DATA5_G12;
  input L_CAM_DATA6_B9;
  input L_CAM_DATA7_A9;
  input L_CAM_DATA8_D9;
  input L_CAM_DATA9_E10;
  input L_CAM_DATA10_B8;
  input L_CAM_DATA11_C7;
  inout  InOut_I2C_L_SDA_B15;
  inout  InOut_I2C_L_SCL_F14;
  inout  InOut_I2C_R_SDA_G9;
  inout  InOut_I2C_R_SCL_F7;


endmodule
